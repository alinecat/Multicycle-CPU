module constant #(parameter V=4, parameter W=32) (out);
	
	output logic [W-1:0]out;
	
	assign out = V ;

endmodule
	