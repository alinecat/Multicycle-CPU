module const_arm #(parameter V=4,W=32) (out);
	
	output logic [W-1:0]out;
	
	assign out = V ;

endmodule
	